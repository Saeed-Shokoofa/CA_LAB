
    



endmodule