module IF(input clk,rst,freeze,Branch_taken, input[31:0] Branch_Addr,output reg [31:0] PC,output [31:0]Instruction );
	reg [7:0]mem[0:128];
	always @(posedge clk, posedge rst)begin
		if(rst) begin
		PC<= 32'b0;
	   ///////////////////////////////////////
	 {mem[0], mem[1], mem[2],    mem[3]}= 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV R0 ,#20 //R0 = 20
     {mem[4], mem[5], mem[6],    mem[7]}= 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV R1 ,#4096 //R1 = 4096
     {mem[8], mem[9], mem[10],    mem[11]}= 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
     {mem[12], mem[13], mem[14],    mem[15]}= 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648
     {mem[16], mem[17], mem[18],    mem[19]}= 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC R4 ,R0,R0 //R4 = 41
     {mem[20], mem[21], mem[22],    mem[23]}= 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
     {mem[24], mem[25], mem[26],    mem[27]}= 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = 10
     {mem[28], mem[29], mem[30],    mem[31]}= 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
     {mem[32], mem[33], mem[34],    mem[35]}= 32'b1110_00_0_0000_0_0111_1000_000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
     {mem[36], mem[37], mem[38],    mem[39]}= 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN R9 ,R6 //R9 = -11
     {mem[40], mem[41], mem[42],    mem[43]}= 32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR R10,R4,R5 //R10 = -84
     {mem[44], mem[45], mem[46],    mem[47]}= 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP R8 ,R6
     {mem[48], mem[49], mem[50],    mem[51]}= 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
     {mem[52], mem[53], mem[54],    mem[55]}= 32'b1110_00_0_1000_1_1001_0000_000000001000; //TST R9 ,R8
     {mem[56], mem[57], mem[58],    mem[59]}= 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
     {mem[60], mem[61], mem[62],    mem[63]}= 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV R0 ,#1024 //R0 = 1024
     {mem[64], mem[65], mem[66],    mem[67]}= 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
     {mem[68], mem[69], mem[70],    mem[71]}= 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR R11,[R0],#0 //R11 = 8192
     {mem[72], mem[73], mem[74],    mem[75]}= 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
     {mem[76], mem[77], mem[78],    mem[79]}= 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
     {mem[80], mem[81], mem[82],    mem[83]}= 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR R4 ,[R0],#13 //MEM[1036] = 41
     {mem[84], mem[85], mem[86],    mem[87]}= 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
     {mem[88], mem[89], mem[90],    mem[91]}= 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
     {mem[92], mem[93], mem[94],    mem[95]}= 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
     {mem[96], mem[97], mem[98],    mem[99]}= 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
     {mem[100], mem[101], mem[102],    mem[103]}= 32'b1110_00_1_1101_0_0000_0001_000000000100; //MOV R1 ,#4 //R1 = 4
     {mem[104], mem[105], mem[106],    mem[107]}= 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV R2 ,#0 //R2 = 0
     {mem[108], mem[109], mem[110],    mem[111]}= 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV R3 ,#0 //R3 = 0
     {mem[112], mem[113], mem[114],    mem[115]}= 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD R4 ,R0,R3,LSL #2
     {mem[116], mem[117], mem[118],    mem[119]}= 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR R5 ,[R4],#0
     {mem[120], mem[121], mem[122],    mem[123]}= 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR R6 ,[R4],#4
     {mem[124], mem[125], mem[126],    mem[127]}= 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP R5 ,R6
     {mem[128], mem[129], mem[130],    mem[131]}= 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT R6 ,[R4],#0
     {mem[132], mem[133], mem[134],    mem[135]}= 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT R5 ,[R4],#4
     {mem[136], mem[137], mem[138],    mem[139]}= 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD R3 ,R3,#1
     {mem[140], mem[141], mem[142],    mem[143]}= 32'b1110_00_1_1010_1_0011_0000_000000000011; //CMP R3 ,#3
     {mem[144], mem[145], mem[146],    mem[147]}= 32'b1011_10_1_0_111111111111111111110111 ; //BLT #-9
     {mem[148], mem[149], mem[150],    mem[151]}= 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD R2 ,R2,#1
     {mem[152], mem[153], mem[154],    mem[155]}= 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP R2 ,R1
     {mem[156], mem[157], mem[158],    mem[159]}= 32'b1011_10_1_0_111111111111111111110011 ; //BLT #-13
     {mem[160], mem[161], mem[162],    mem[163]}= 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
     {mem[164], mem[165], mem[166],    mem[167]}= 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
     {mem[168], mem[169], mem[170],    mem[171]}= 32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR R3 ,[R0],#8 //R3 = 41
	 {mem[172], mem[173], mem[174],    mem[175]}= 32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR R4 ,[R0],#12 //R4 = 8192
     {mem[176], mem[177], mem[178],    mem[179]}= 32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR R5 ,[R0],#16 //R5 = -123
     {mem[180], mem[181], mem[182],    mem[183]}= 32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR R6 ,[R0],#20 //R4 = 10
     {mem[184], mem[185], mem[186],    mem[187]}= 32'b1110_10_1_0_111111111111111111111111 ; //B #-1
	   ///////////////////////////////////////
	 end
		else begin
			PC<=PC+32'd4;
		end
	end
	assign Instruction = {mem[PC], mem[PC+32'd1], mem[PC+32'd2], mem[PC+32'd3]};
endmodule
