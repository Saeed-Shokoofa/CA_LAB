module ARM(clk,rst);

input clk,rst;
wire if_br_taken,exe_br_taken,id_z,id_c,id_n,id_v,id_WB_EN,id_MEM_R,id_MEM_W,id_B,id_S,id_imm
wire [3:0]id_EXE_CMD,id_dest
wire [11:0]id_shift_operand;
wire [23:0]id_signed_imm
wire[31:0]if_br_adr,if_pc,if_inst,if_pc_out,if_inst_out,id_PC,id_val_rn,id_val_rm,


IF IF_stg(.clk(clk),.rst(rst),.freeze(1'b0),.Branch_taken(if_br_taken),.Branch_Addr(if_br_adr),.PC(if_pc),.Instruction(if_inst));
IF_reg IF_register(.clk(clk),.rst(rst),.freeze(1'b0),.flush(exe_br_taken),.PC_in(if_pc),.Instruction_in(if_inst),.PC(if_pc_out),.Instruction(if_inst_out));
ID ID_stg(.clk(clk),.rst(rst),.z(id_z),.c(id_c),.n(id_n),.v(id_v),.instruction(if_inst_out),.PC(if_pc_out),.WB_WB_EN(),.WB_Value(),.WB_Dest(),.
    WB_EN(id_WB_EN),.MEM_R(id_MEM_R),.MEM_W(id_MEM_W),.EXE_CMD(id_EXE_CMD),.B(id_B),.S(id_S),.PC_out(id_PC),.val_rn(id_val_rn),.val_rm(id_val_rm),.dest(id_dest),.signed_imm(id_signed_imm),.imm(id_imm),.Shift_Operand(id_shift_operand));
ID_REG ID_rsgister(.clk(clk),.rst(rst),.flush(exe_br_taken),.carry(),.dest(),.signed_imm(),.Shift_Operand(),.imm(),.val_rm(),.val_rn(),.PC(),.S(),.B(),.EXE_CMD(),.MEM_W(),.MEM_R(),.WB_EN(),.
    carry_out(),.dest_out(),.signed_imm_out(),.Shift_Operand_out(),.imm_out(),.val_rm_out(),.val_rn_out(),.PC_out(),.S_out(),.B_out(),.
    EXE_CMD_out(),.MEM_W_out(),.MEM_R_out(),.WB_EN_out());
EXE EXE_stg(.clk(clk),.rst(rst),.WB_EN(),.MEM_R(),.MEM_W(),.EXE_CMD(),.B(),.S(),.PC(),.val_rn(),.val_rm(),.imm(),.Shift_Operand(),.signed_imm(),.dest(),.carry(),.
    WB_EN_out(),.MEM_R_out(),.MEM_W_out(),.ALU_res(),.val_rm_out(),.dest_out(),.branch_adr(),.status_out(),.branch_taken(exe_br_taken));
EXE_reg EXE_register(.clk(clk),.rst(rst),.dest(),.val_rm(),.ALU_res(),.MEM_W(),.MEM_R(),.WB_EN(),.
    dest_out(),.val_rm_out(),.ALU_res_out(),.MEM_W_out(),.MEM_R_out(),.WB_EN_out());

endmodule